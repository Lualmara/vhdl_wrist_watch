----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 18.11.2021 01:16:40
-- Design Name: 
-- Module Name: wristwatch_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity wristwatch_tb is
--  Port ( );
end wristwatch_tb;

architecture Behavioral of wristwatch_tb is

component main is
    PORT(

		mode : in STD_LOGIC;
		config : in STD_LOGIC_VECTOR(1 DOWNTO 0);
		chv0 : in STD_LOGIC; -- por enquanto nao faz nada
		
		chrono_start : in STD_LOGIC;
		chrono_stop : in STD_LOGIC;
		chrono_reset : in STD_LOGIC;
		
		seg_unid : OUT STD_LOGIC_VECTOR(6 downto 0);
		seg_dez : OUT STD_LOGIC_VECTOR(6 downto 0);
		min_unid : OUT STD_LOGIC_VECTOR(6 downto 0);
		min_dez : OUT STD_LOGIC_VECTOR(6 downto 0);
		hora_unid : OUT STD_LOGIC_VECTOR(6 downto 0);
		hora_dez : OUT STD_LOGIC_VECTOR(6 downto 0);
		am_pm : OUT STD_LOGIC;

	);
end component;

constant clk;
signal mode, config, chv0, chrono_start, chrono_stop, chrono_reset, ;

begin


end Behavioral;
